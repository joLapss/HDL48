-- lab2q.vhd

-- Generated using ACDS version 14.1 186 at 2015.05.24.13:51:31

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lab2q is
	port (
		clk_clk       : in    std_logic                     := '0';             --       clk.clk
		clk_sdram_clk : out   std_logic;                                        -- clk_sdram.clk
		mouse_CLK     : inout std_logic                     := '0';             --     mouse.CLK
		mouse_DAT     : inout std_logic                     := '0';             --          .DAT
		reset_reset_n : in    std_logic                     := '0';             --     reset.reset_n
		sram_addr     : out   std_logic_vector(12 downto 0);                    --      sram.addr
		sram_ba       : out   std_logic_vector(1 downto 0);                     --          .ba
		sram_cas_n    : out   std_logic;                                        --          .cas_n
		sram_cke      : out   std_logic;                                        --          .cke
		sram_cs_n     : out   std_logic;                                        --          .cs_n
		sram_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sram_dqm      : out   std_logic_vector(1 downto 0);                     --          .dqm
		sram_ras_n    : out   std_logic;                                        --          .ras_n
		sram_we_n     : out   std_logic;                                        --          .we_n
		vga_out_CLK   : out   std_logic;                                        --   vga_out.CLK
		vga_out_HS    : out   std_logic;                                        --          .HS
		vga_out_VS    : out   std_logic;                                        --          .VS
		vga_out_BLANK : out   std_logic;                                        --          .BLANK
		vga_out_SYNC  : out   std_logic;                                        --          .SYNC
		vga_out_R     : out   std_logic_vector(7 downto 0);                     --          .R
		vga_out_G     : out   std_logic_vector(7 downto 0);                     --          .G
		vga_out_B     : out   std_logic_vector(7 downto 0)                      --          .B
	);
end entity lab2q;

architecture rtl of lab2q is
	component lab2q_blender is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			foreground_data          : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			foreground_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			foreground_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			foreground_valid         : in  std_logic                     := 'X';             -- valid
			foreground_ready         : out std_logic;                                        -- ready
			background_data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			background_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			background_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			background_valid         : in  std_logic                     := 'X';             -- valid
			background_ready         : out std_logic;                                        -- ready
			output_ready             : in  std_logic                     := 'X';             -- ready
			output_data              : out std_logic_vector(29 downto 0);                    -- data
			output_startofpacket     : out std_logic;                                        -- startofpacket
			output_endofpacket       : out std_logic;                                        -- endofpacket
			output_valid             : out std_logic                                         -- valid
		);
	end component lab2q_blender;

	component lab2q_character_buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(39 downto 0)                     -- data
		);
	end component lab2q_character_buffer;

	component lab2q_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component lab2q_cpu;

	component lab2q_fifo is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component lab2q_fifo;

	component lab2q_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component lab2q_jtag_uart;

	component lab2q_mouse_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component lab2q_mouse_0;

	component lab2q_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component lab2q_onchip_mem;

	component lab2q_pixel_buffer is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component lab2q_pixel_buffer;

	component lab2q_resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component lab2q_resampler;

	component lab2q_scaler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component lab2q_scaler;

	component lab2q_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component lab2q_sdram_controller;

	component lab2q_sys_sdram_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component lab2q_sys_sdram_pll;

	component lab2q_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component lab2q_sysid;

	component lab2q_vga_controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component lab2q_vga_controller;

	component lab2q_video_clk is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			video_in_clk_clk   : out std_logic;        -- clk
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component lab2q_video_clk;

	component lab2q_mm_interconnect_0 is
		port (
			sys_sdram_pll_sys_clk_clk                          : in  std_logic                     := 'X';             -- clk
			pixel_buffer_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			pixel_buffer_avalon_pixel_dma_master_address       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			pixel_buffer_avalon_pixel_dma_master_waitrequest   : out std_logic;                                        -- waitrequest
			pixel_buffer_avalon_pixel_dma_master_read          : in  std_logic                     := 'X';             -- read
			pixel_buffer_avalon_pixel_dma_master_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			pixel_buffer_avalon_pixel_dma_master_readdatavalid : out std_logic;                                        -- readdatavalid
			pixel_buffer_avalon_pixel_dma_master_lock          : in  std_logic                     := 'X';             -- lock
			onchip_mem_s1_address                              : out std_logic_vector(15 downto 0);                    -- address
			onchip_mem_s1_write                                : out std_logic;                                        -- write
			onchip_mem_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                           : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                                : out std_logic                                         -- clken
		);
	end component lab2q_mm_interconnect_0;

	component lab2q_mm_interconnect_1 is
		port (
			sys_sdram_pll_sys_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			sysid_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                  : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                 : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			character_buffer_avalon_char_buffer_slave_address     : out std_logic_vector(12 downto 0);                    -- address
			character_buffer_avalon_char_buffer_slave_write       : out std_logic;                                        -- write
			character_buffer_avalon_char_buffer_slave_read        : out std_logic;                                        -- read
			character_buffer_avalon_char_buffer_slave_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			character_buffer_avalon_char_buffer_slave_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			character_buffer_avalon_char_buffer_slave_byteenable  : out std_logic_vector(0 downto 0);                     -- byteenable
			character_buffer_avalon_char_buffer_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			character_buffer_avalon_char_buffer_slave_chipselect  : out std_logic;                                        -- chipselect
			character_buffer_avalon_char_control_slave_address    : out std_logic_vector(0 downto 0);                     -- address
			character_buffer_avalon_char_control_slave_write      : out std_logic;                                        -- write
			character_buffer_avalon_char_control_slave_read       : out std_logic;                                        -- read
			character_buffer_avalon_char_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			character_buffer_avalon_char_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			character_buffer_avalon_char_control_slave_byteenable : out std_logic_vector(3 downto 0);                     -- byteenable
			character_buffer_avalon_char_control_slave_chipselect : out std_logic;                                        -- chipselect
			cpu_jtag_debug_module_address                         : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write                           : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                            : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess                     : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			mouse_0_avalon_ps2_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			mouse_0_avalon_ps2_slave_write                        : out std_logic;                                        -- write
			mouse_0_avalon_ps2_slave_read                         : out std_logic;                                        -- read
			mouse_0_avalon_ps2_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mouse_0_avalon_ps2_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			mouse_0_avalon_ps2_slave_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			mouse_0_avalon_ps2_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			mouse_0_avalon_ps2_slave_chipselect                   : out std_logic;                                        -- chipselect
			pixel_buffer_avalon_control_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			pixel_buffer_avalon_control_slave_write               : out std_logic;                                        -- write
			pixel_buffer_avalon_control_slave_read                : out std_logic;                                        -- read
			pixel_buffer_avalon_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pixel_buffer_avalon_control_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			pixel_buffer_avalon_control_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_controller_s1_address                           : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                             : out std_logic;                                        -- write
			sdram_controller_s1_read                              : out std_logic;                                        -- read
			sdram_controller_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                        : out std_logic;                                        -- chipselect
			sysid_control_slave_address                           : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component lab2q_mm_interconnect_1;

	component lab2q_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component lab2q_irq_mapper;

	component lab2q_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component lab2q_rst_controller;

	component lab2q_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component lab2q_rst_controller_001;

	signal blender_avalon_blended_source_valid                                     : std_logic;                     -- blender:output_valid -> fifo:stream_in_valid
	signal blender_avalon_blended_source_data                                      : std_logic_vector(29 downto 0); -- blender:output_data -> fifo:stream_in_data
	signal blender_avalon_blended_source_ready                                     : std_logic;                     -- fifo:stream_in_ready -> blender:output_ready
	signal blender_avalon_blended_source_startofpacket                             : std_logic;                     -- blender:output_startofpacket -> fifo:stream_in_startofpacket
	signal blender_avalon_blended_source_endofpacket                               : std_logic;                     -- blender:output_endofpacket -> fifo:stream_in_endofpacket
	signal character_buffer_avalon_char_source_valid                               : std_logic;                     -- character_buffer:stream_valid -> blender:foreground_valid
	signal character_buffer_avalon_char_source_data                                : std_logic_vector(39 downto 0); -- character_buffer:stream_data -> blender:foreground_data
	signal character_buffer_avalon_char_source_ready                               : std_logic;                     -- blender:foreground_ready -> character_buffer:stream_ready
	signal character_buffer_avalon_char_source_startofpacket                       : std_logic;                     -- character_buffer:stream_startofpacket -> blender:foreground_startofpacket
	signal character_buffer_avalon_char_source_endofpacket                         : std_logic;                     -- character_buffer:stream_endofpacket -> blender:foreground_endofpacket
	signal fifo_avalon_dc_buffer_source_valid                                      : std_logic;                     -- fifo:stream_out_valid -> vga_controller:valid
	signal fifo_avalon_dc_buffer_source_data                                       : std_logic_vector(29 downto 0); -- fifo:stream_out_data -> vga_controller:data
	signal fifo_avalon_dc_buffer_source_ready                                      : std_logic;                     -- vga_controller:ready -> fifo:stream_out_ready
	signal fifo_avalon_dc_buffer_source_startofpacket                              : std_logic;                     -- fifo:stream_out_startofpacket -> vga_controller:startofpacket
	signal fifo_avalon_dc_buffer_source_endofpacket                                : std_logic;                     -- fifo:stream_out_endofpacket -> vga_controller:endofpacket
	signal pixel_buffer_avalon_pixel_source_valid                                  : std_logic;                     -- pixel_buffer:stream_valid -> resampler:stream_in_valid
	signal pixel_buffer_avalon_pixel_source_data                                   : std_logic_vector(15 downto 0); -- pixel_buffer:stream_data -> resampler:stream_in_data
	signal pixel_buffer_avalon_pixel_source_ready                                  : std_logic;                     -- resampler:stream_in_ready -> pixel_buffer:stream_ready
	signal pixel_buffer_avalon_pixel_source_startofpacket                          : std_logic;                     -- pixel_buffer:stream_startofpacket -> resampler:stream_in_startofpacket
	signal pixel_buffer_avalon_pixel_source_endofpacket                            : std_logic;                     -- pixel_buffer:stream_endofpacket -> resampler:stream_in_endofpacket
	signal resampler_avalon_rgb_source_valid                                       : std_logic;                     -- resampler:stream_out_valid -> scaler:stream_in_valid
	signal resampler_avalon_rgb_source_data                                        : std_logic_vector(29 downto 0); -- resampler:stream_out_data -> scaler:stream_in_data
	signal resampler_avalon_rgb_source_ready                                       : std_logic;                     -- scaler:stream_in_ready -> resampler:stream_out_ready
	signal resampler_avalon_rgb_source_startofpacket                               : std_logic;                     -- resampler:stream_out_startofpacket -> scaler:stream_in_startofpacket
	signal resampler_avalon_rgb_source_endofpacket                                 : std_logic;                     -- resampler:stream_out_endofpacket -> scaler:stream_in_endofpacket
	signal scaler_avalon_scaler_source_valid                                       : std_logic;                     -- scaler:stream_out_valid -> blender:background_valid
	signal scaler_avalon_scaler_source_data                                        : std_logic_vector(29 downto 0); -- scaler:stream_out_data -> blender:background_data
	signal scaler_avalon_scaler_source_ready                                       : std_logic;                     -- blender:background_ready -> scaler:stream_out_ready
	signal scaler_avalon_scaler_source_startofpacket                               : std_logic;                     -- scaler:stream_out_startofpacket -> blender:background_startofpacket
	signal scaler_avalon_scaler_source_endofpacket                                 : std_logic;                     -- scaler:stream_out_endofpacket -> blender:background_endofpacket
	signal sys_sdram_pll_sys_clk_clk                                               : std_logic;                     -- sys_sdram_pll:sys_clk_clk -> [blender:clk, character_buffer:clk, cpu:clk, fifo:clk_stream_in, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:sys_sdram_pll_sys_clk_clk, mm_interconnect_1:sys_sdram_pll_sys_clk_clk, mouse_0:clk, onchip_mem:clk, pixel_buffer:clk, resampler:clk, rst_controller:clk, rst_controller_002:clk, scaler:clk, sdram_controller:clk, sysid:clock]
	signal video_clk_vga_clk_clk                                                   : std_logic;                     -- video_clk:vga_clk_clk -> [fifo:clk_stream_out, rst_controller_001:clk, vga_controller:clk]
	signal pixel_buffer_avalon_pixel_dma_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_waitrequest -> pixel_buffer:master_waitrequest
	signal pixel_buffer_avalon_pixel_dma_master_readdata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_readdata -> pixel_buffer:master_readdata
	signal pixel_buffer_avalon_pixel_dma_master_address                            : std_logic_vector(31 downto 0); -- pixel_buffer:master_address -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_address
	signal pixel_buffer_avalon_pixel_dma_master_read                               : std_logic;                     -- pixel_buffer:master_read -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_read
	signal pixel_buffer_avalon_pixel_dma_master_readdatavalid                      : std_logic;                     -- mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_readdatavalid -> pixel_buffer:master_readdatavalid
	signal pixel_buffer_avalon_pixel_dma_master_lock                               : std_logic;                     -- pixel_buffer:master_arbiterlock -> mm_interconnect_0:pixel_buffer_avalon_pixel_dma_master_lock
	signal mm_interconnect_0_onchip_mem_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                                : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                                   : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                                   : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal cpu_data_master_readdata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                             : std_logic;                     -- mm_interconnect_1:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                             : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_1:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                 : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_1:cpu_data_master_address
	signal cpu_data_master_byteenable                                              : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_1:cpu_data_master_byteenable
	signal cpu_data_master_read                                                    : std_logic;                     -- cpu:d_read -> mm_interconnect_1:cpu_data_master_read
	signal cpu_data_master_write                                                   : std_logic;                     -- cpu:d_write -> mm_interconnect_1:cpu_data_master_write
	signal cpu_data_master_writedata                                               : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_1:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                      : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                          : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	signal cpu_instruction_master_read                                             : std_logic;                     -- cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                    : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_chipselect  : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_chipselect -> character_buffer:buf_chipselect
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_readdata    : std_logic_vector(7 downto 0);  -- character_buffer:buf_readdata -> mm_interconnect_1:character_buffer_avalon_char_buffer_slave_readdata
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_waitrequest : std_logic;                     -- character_buffer:buf_waitrequest -> mm_interconnect_1:character_buffer_avalon_char_buffer_slave_waitrequest
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_address     : std_logic_vector(12 downto 0); -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_address -> character_buffer:buf_address
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_read        : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_read -> character_buffer:buf_read
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_byteenable  : std_logic_vector(0 downto 0);  -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_byteenable -> character_buffer:buf_byteenable
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_write       : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_write -> character_buffer:buf_write
	signal mm_interconnect_1_character_buffer_avalon_char_buffer_slave_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_1:character_buffer_avalon_char_buffer_slave_writedata -> character_buffer:buf_writedata
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_chipselect : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_control_slave_chipselect -> character_buffer:ctrl_chipselect
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_readdata   : std_logic_vector(31 downto 0); -- character_buffer:ctrl_readdata -> mm_interconnect_1:character_buffer_avalon_char_control_slave_readdata
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_address    : std_logic_vector(0 downto 0);  -- mm_interconnect_1:character_buffer_avalon_char_control_slave_address -> character_buffer:ctrl_address
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_read       : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_control_slave_read -> character_buffer:ctrl_read
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_1:character_buffer_avalon_char_control_slave_byteenable -> character_buffer:ctrl_byteenable
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_write      : std_logic;                     -- mm_interconnect_1:character_buffer_avalon_char_control_slave_write -> character_buffer:ctrl_write
	signal mm_interconnect_1_character_buffer_avalon_char_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_1:character_buffer_avalon_char_control_slave_writedata -> character_buffer:ctrl_writedata
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_readdata            : std_logic_vector(31 downto 0); -- pixel_buffer:slave_readdata -> mm_interconnect_1:pixel_buffer_avalon_control_slave_readdata
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_1:pixel_buffer_avalon_control_slave_address -> pixel_buffer:slave_address
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_read                : std_logic;                     -- mm_interconnect_1:pixel_buffer_avalon_control_slave_read -> pixel_buffer:slave_read
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_1:pixel_buffer_avalon_control_slave_byteenable -> pixel_buffer:slave_byteenable
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_write               : std_logic;                     -- mm_interconnect_1:pixel_buffer_avalon_control_slave_write -> pixel_buffer:slave_write
	signal mm_interconnect_1_pixel_buffer_avalon_control_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_1:pixel_buffer_avalon_control_slave_writedata -> pixel_buffer:slave_writedata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect                : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata                  : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest               : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read                      : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write                     : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_chipselect                   : std_logic;                     -- mm_interconnect_1:mouse_0_avalon_ps2_slave_chipselect -> mouse_0:chipselect
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_readdata                     : std_logic_vector(31 downto 0); -- mouse_0:readdata -> mm_interconnect_1:mouse_0_avalon_ps2_slave_readdata
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_waitrequest                  : std_logic;                     -- mouse_0:waitrequest -> mm_interconnect_1:mouse_0_avalon_ps2_slave_waitrequest
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_1:mouse_0_avalon_ps2_slave_address -> mouse_0:address
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_read                         : std_logic;                     -- mm_interconnect_1:mouse_0_avalon_ps2_slave_read -> mouse_0:read
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:mouse_0_avalon_ps2_slave_byteenable -> mouse_0:byteenable
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_write                        : std_logic;                     -- mm_interconnect_1:mouse_0_avalon_ps2_slave_write -> mouse_0:write
	signal mm_interconnect_1_mouse_0_avalon_ps2_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:mouse_0_avalon_ps2_slave_writedata -> mouse_0:writedata
	signal mm_interconnect_1_sysid_control_slave_readdata                          : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	signal mm_interconnect_1_sysid_control_slave_address                           : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_1_cpu_jtag_debug_module_readdata                        : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_1:cpu_jtag_debug_module_readdata
	signal mm_interconnect_1_cpu_jtag_debug_module_waitrequest                     : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_1:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_1_cpu_jtag_debug_module_debugaccess                     : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_1_cpu_jtag_debug_module_address                         : std_logic_vector(8 downto 0);  -- mm_interconnect_1:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_1_cpu_jtag_debug_module_read                            : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_1_cpu_jtag_debug_module_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_1:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_1_cpu_jtag_debug_module_write                           : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_1_cpu_jtag_debug_module_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_1_sdram_controller_s1_chipselect                        : std_logic;                     -- mm_interconnect_1:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_1_sdram_controller_s1_readdata                          : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_1:sdram_controller_s1_readdata
	signal mm_interconnect_1_sdram_controller_s1_waitrequest                       : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_1:sdram_controller_s1_waitrequest
	signal mm_interconnect_1_sdram_controller_s1_address                           : std_logic_vector(24 downto 0); -- mm_interconnect_1:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_1_sdram_controller_s1_read                              : std_logic;                     -- mm_interconnect_1:sdram_controller_s1_read -> mm_interconnect_1_sdram_controller_s1_read:in
	signal mm_interconnect_1_sdram_controller_s1_byteenable                        : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sdram_controller_s1_byteenable -> mm_interconnect_1_sdram_controller_s1_byteenable:in
	signal mm_interconnect_1_sdram_controller_s1_readdatavalid                     : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_1:sdram_controller_s1_readdatavalid
	signal mm_interconnect_1_sdram_controller_s1_write                             : std_logic;                     -- mm_interconnect_1:sdram_controller_s1_write -> mm_interconnect_1_sdram_controller_s1_write:in
	signal mm_interconnect_1_sdram_controller_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_1:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal irq_mapper_receiver0_irq                                                : std_logic;                     -- mouse_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal rst_controller_reset_out_reset                                          : std_logic;                     -- rst_controller:reset_out -> [blender:reset, character_buffer:reset, fifo:reset_stream_in, irq_mapper:reset, mm_interconnect_0:pixel_buffer_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_n_reset_bridge_in_reset_reset, mouse_0:reset, onchip_mem:reset, pixel_buffer:reset, resampler:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, scaler:reset]
	signal rst_controller_reset_out_reset_req                                      : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal sys_sdram_pll_reset_source_reset                                        : std_logic;                     -- sys_sdram_pll:reset_source_reset -> rst_controller:reset_in0
	signal rst_controller_001_reset_out_reset                                      : std_logic;                     -- rst_controller_001:reset_out -> [fifo:reset_stream_out, vga_controller:reset]
	signal video_clk_reset_source_reset                                            : std_logic;                     -- video_clk:reset_source_reset -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                                      : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_1:sysid_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                                 : std_logic;                     -- reset_reset_n:inv -> [rst_controller_002:reset_in0, sys_sdram_pll:ref_reset_reset, video_clk:ref_reset_reset]
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv            : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv           : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_1_sdram_controller_s1_read_ports_inv                    : std_logic;                     -- mm_interconnect_1_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_1_sdram_controller_s1_byteenable_ports_inv              : std_logic_vector(1 downto 0);  -- mm_interconnect_1_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_1_sdram_controller_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_1_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n]
	signal rst_controller_002_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [sdram_controller:reset_n, sysid:reset_n]

begin

	blender : component lab2q_blender
		port map (
			clk                      => sys_sdram_pll_sys_clk_clk,                         --                    clk.clk
			reset                    => rst_controller_reset_out_reset,                    --                  reset.reset
			foreground_data          => character_buffer_avalon_char_source_data,          -- avalon_foreground_sink.data
			foreground_startofpacket => character_buffer_avalon_char_source_startofpacket, --                       .startofpacket
			foreground_endofpacket   => character_buffer_avalon_char_source_endofpacket,   --                       .endofpacket
			foreground_valid         => character_buffer_avalon_char_source_valid,         --                       .valid
			foreground_ready         => character_buffer_avalon_char_source_ready,         --                       .ready
			background_data          => scaler_avalon_scaler_source_data,                  -- avalon_background_sink.data
			background_startofpacket => scaler_avalon_scaler_source_startofpacket,         --                       .startofpacket
			background_endofpacket   => scaler_avalon_scaler_source_endofpacket,           --                       .endofpacket
			background_valid         => scaler_avalon_scaler_source_valid,                 --                       .valid
			background_ready         => scaler_avalon_scaler_source_ready,                 --                       .ready
			output_ready             => blender_avalon_blended_source_ready,               --  avalon_blended_source.ready
			output_data              => blender_avalon_blended_source_data,                --                       .data
			output_startofpacket     => blender_avalon_blended_source_startofpacket,       --                       .startofpacket
			output_endofpacket       => blender_avalon_blended_source_endofpacket,         --                       .endofpacket
			output_valid             => blender_avalon_blended_source_valid                --                       .valid
		);

	character_buffer : component lab2q_character_buffer
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                                 --                       clk.clk
			reset                => rst_controller_reset_out_reset,                                            --                     reset.reset
			ctrl_address         => mm_interconnect_1_character_buffer_avalon_char_control_slave_address(0),   -- avalon_char_control_slave.address
			ctrl_byteenable      => mm_interconnect_1_character_buffer_avalon_char_control_slave_byteenable,   --                          .byteenable
			ctrl_chipselect      => mm_interconnect_1_character_buffer_avalon_char_control_slave_chipselect,   --                          .chipselect
			ctrl_read            => mm_interconnect_1_character_buffer_avalon_char_control_slave_read,         --                          .read
			ctrl_write           => mm_interconnect_1_character_buffer_avalon_char_control_slave_write,        --                          .write
			ctrl_writedata       => mm_interconnect_1_character_buffer_avalon_char_control_slave_writedata,    --                          .writedata
			ctrl_readdata        => mm_interconnect_1_character_buffer_avalon_char_control_slave_readdata,     --                          .readdata
			buf_byteenable       => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_byteenable(0), --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_chipselect,    --                          .chipselect
			buf_read             => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_read,          --                          .read
			buf_write            => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_write,         --                          .write
			buf_writedata        => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_writedata,     --                          .writedata
			buf_readdata         => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_readdata,      --                          .readdata
			buf_waitrequest      => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_waitrequest,   --                          .waitrequest
			buf_address          => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_address,       --                          .address
			stream_ready         => character_buffer_avalon_char_source_ready,                                 --        avalon_char_source.ready
			stream_startofpacket => character_buffer_avalon_char_source_startofpacket,                         --                          .startofpacket
			stream_endofpacket   => character_buffer_avalon_char_source_endofpacket,                           --                          .endofpacket
			stream_valid         => character_buffer_avalon_char_source_valid,                                 --                          .valid
			stream_data          => character_buffer_avalon_char_source_data                                   --                          .data
		);

	cpu : component lab2q_cpu
		port map (
			clk                                   => sys_sdram_pll_sys_clk_clk,                           --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_1_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_1_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_1_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_1_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_1_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_1_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_1_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_1_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	fifo : component lab2q_fifo
		port map (
			clk_stream_in            => sys_sdram_pll_sys_clk_clk,                   --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,              --         reset_stream_in.reset
			clk_stream_out           => video_clk_vga_clk_clk,                       --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,          --        reset_stream_out.reset
			stream_in_ready          => blender_avalon_blended_source_ready,         --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => blender_avalon_blended_source_startofpacket, --                        .startofpacket
			stream_in_endofpacket    => blender_avalon_blended_source_endofpacket,   --                        .endofpacket
			stream_in_valid          => blender_avalon_blended_source_valid,         --                        .valid
			stream_in_data           => blender_avalon_blended_source_data,          --                        .data
			stream_out_ready         => fifo_avalon_dc_buffer_source_ready,          -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => fifo_avalon_dc_buffer_source_startofpacket,  --                        .startofpacket
			stream_out_endofpacket   => fifo_avalon_dc_buffer_source_endofpacket,    --                        .endofpacket
			stream_out_valid         => fifo_avalon_dc_buffer_source_valid,          --                        .valid
			stream_out_data          => fifo_avalon_dc_buffer_source_data            --                        .data
		);

	jtag_uart : component lab2q_jtag_uart
		port map (
			clk            => sys_sdram_pll_sys_clk_clk,                                     --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	mouse_0 : component lab2q_mouse_0
		port map (
			clk         => sys_sdram_pll_sys_clk_clk,                              --                clk.clk
			reset       => rst_controller_reset_out_reset,                         --              reset.reset
			address     => mm_interconnect_1_mouse_0_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_1_mouse_0_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_1_mouse_0_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_1_mouse_0_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_1_mouse_0_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_1_mouse_0_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_1_mouse_0_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_1_mouse_0_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => irq_mapper_receiver0_irq,                               --          interrupt.irq
			PS2_CLK     => mouse_CLK,                                              -- external_interface.export
			PS2_DAT     => mouse_DAT                                               --                   .export
		);

	onchip_mem : component lab2q_onchip_mem
		port map (
			clk        => sys_sdram_pll_sys_clk_clk,                  --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	pixel_buffer : component lab2q_pixel_buffer
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                      --                     clk.clk
			reset                => rst_controller_reset_out_reset,                                 --                   reset.reset
			master_readdatavalid => pixel_buffer_avalon_pixel_dma_master_readdatavalid,             -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => pixel_buffer_avalon_pixel_dma_master_waitrequest,               --                        .waitrequest
			master_address       => pixel_buffer_avalon_pixel_dma_master_address,                   --                        .address
			master_arbiterlock   => pixel_buffer_avalon_pixel_dma_master_lock,                      --                        .lock
			master_read          => pixel_buffer_avalon_pixel_dma_master_read,                      --                        .read
			master_readdata      => pixel_buffer_avalon_pixel_dma_master_readdata,                  --                        .readdata
			slave_address        => mm_interconnect_1_pixel_buffer_avalon_control_slave_address,    --    avalon_control_slave.address
			slave_byteenable     => mm_interconnect_1_pixel_buffer_avalon_control_slave_byteenable, --                        .byteenable
			slave_read           => mm_interconnect_1_pixel_buffer_avalon_control_slave_read,       --                        .read
			slave_write          => mm_interconnect_1_pixel_buffer_avalon_control_slave_write,      --                        .write
			slave_writedata      => mm_interconnect_1_pixel_buffer_avalon_control_slave_writedata,  --                        .writedata
			slave_readdata       => mm_interconnect_1_pixel_buffer_avalon_control_slave_readdata,   --                        .readdata
			stream_ready         => pixel_buffer_avalon_pixel_source_ready,                         --     avalon_pixel_source.ready
			stream_startofpacket => pixel_buffer_avalon_pixel_source_startofpacket,                 --                        .startofpacket
			stream_endofpacket   => pixel_buffer_avalon_pixel_source_endofpacket,                   --                        .endofpacket
			stream_valid         => pixel_buffer_avalon_pixel_source_valid,                         --                        .valid
			stream_data          => pixel_buffer_avalon_pixel_source_data                           --                        .data
		);

	resampler : component lab2q_resampler
		port map (
			clk                      => sys_sdram_pll_sys_clk_clk,                      --               clk.clk
			reset                    => rst_controller_reset_out_reset,                 --             reset.reset
			stream_in_startofpacket  => pixel_buffer_avalon_pixel_source_startofpacket, --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => pixel_buffer_avalon_pixel_source_endofpacket,   --                  .endofpacket
			stream_in_valid          => pixel_buffer_avalon_pixel_source_valid,         --                  .valid
			stream_in_ready          => pixel_buffer_avalon_pixel_source_ready,         --                  .ready
			stream_in_data           => pixel_buffer_avalon_pixel_source_data,          --                  .data
			stream_out_ready         => resampler_avalon_rgb_source_ready,              -- avalon_rgb_source.ready
			stream_out_startofpacket => resampler_avalon_rgb_source_startofpacket,      --                  .startofpacket
			stream_out_endofpacket   => resampler_avalon_rgb_source_endofpacket,        --                  .endofpacket
			stream_out_valid         => resampler_avalon_rgb_source_valid,              --                  .valid
			stream_out_data          => resampler_avalon_rgb_source_data                --                  .data
		);

	scaler : component lab2q_scaler
		port map (
			clk                      => sys_sdram_pll_sys_clk_clk,                 --                  clk.clk
			reset                    => rst_controller_reset_out_reset,            --                reset.reset
			stream_in_startofpacket  => resampler_avalon_rgb_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => resampler_avalon_rgb_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => resampler_avalon_rgb_source_valid,         --                     .valid
			stream_in_ready          => resampler_avalon_rgb_source_ready,         --                     .ready
			stream_in_data           => resampler_avalon_rgb_source_data,          --                     .data
			stream_out_ready         => scaler_avalon_scaler_source_ready,         -- avalon_scaler_source.ready
			stream_out_startofpacket => scaler_avalon_scaler_source_startofpacket, --                     .startofpacket
			stream_out_endofpacket   => scaler_avalon_scaler_source_endofpacket,   --                     .endofpacket
			stream_out_valid         => scaler_avalon_scaler_source_valid,         --                     .valid
			stream_out_data          => scaler_avalon_scaler_source_data           --                     .data
		);

	sdram_controller : component lab2q_sdram_controller
		port map (
			clk            => sys_sdram_pll_sys_clk_clk,                                  --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,               -- reset.reset_n
			az_addr        => mm_interconnect_1_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_1_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_1_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_1_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_1_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_1_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_1_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_1_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_1_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sram_addr,                                                  --  wire.export
			zs_ba          => sram_ba,                                                    --      .export
			zs_cas_n       => sram_cas_n,                                                 --      .export
			zs_cke         => sram_cke,                                                   --      .export
			zs_cs_n        => sram_cs_n,                                                  --      .export
			zs_dq          => sram_dq,                                                    --      .export
			zs_dqm         => sram_dqm,                                                   --      .export
			zs_ras_n       => sram_ras_n,                                                 --      .export
			zs_we_n        => sram_we_n                                                   --      .export
		);

	sys_sdram_pll : component lab2q_sys_sdram_pll
		port map (
			ref_clk_clk        => clk_clk,                          --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,          --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => clk_sdram_clk,                    --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_reset_source_reset  -- reset_source.reset
		);

	sysid : component lab2q_sysid
		port map (
			clock    => sys_sdram_pll_sys_clk_clk,                        --           clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_1_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_control_slave_address(0)  --              .address
		);

	vga_controller : component lab2q_vga_controller
		port map (
			clk           => video_clk_vga_clk_clk,                      --                clk.clk
			reset         => rst_controller_001_reset_out_reset,         --              reset.reset
			data          => fifo_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => fifo_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => fifo_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => fifo_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => fifo_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_out_CLK,                                -- external_interface.export
			VGA_HS        => vga_out_HS,                                 --                   .export
			VGA_VS        => vga_out_VS,                                 --                   .export
			VGA_BLANK     => vga_out_BLANK,                              --                   .export
			VGA_SYNC      => vga_out_SYNC,                               --                   .export
			VGA_R         => vga_out_R,                                  --                   .export
			VGA_G         => vga_out_G,                                  --                   .export
			VGA_B         => vga_out_B                                   --                   .export
		);

	video_clk : component lab2q_video_clk
		port map (
			ref_clk_clk        => clk_clk,                      --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,      --    ref_reset.reset
			video_in_clk_clk   => open,                         -- video_in_clk.clk
			vga_clk_clk        => video_clk_vga_clk_clk,        --      vga_clk.clk
			reset_source_reset => video_clk_reset_source_reset  -- reset_source.reset
		);

	mm_interconnect_0 : component lab2q_mm_interconnect_0
		port map (
			sys_sdram_pll_sys_clk_clk                          => sys_sdram_pll_sys_clk_clk,                          --                    sys_sdram_pll_sys_clk.clk
			pixel_buffer_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                     -- pixel_buffer_reset_reset_bridge_in_reset.reset
			pixel_buffer_avalon_pixel_dma_master_address       => pixel_buffer_avalon_pixel_dma_master_address,       --     pixel_buffer_avalon_pixel_dma_master.address
			pixel_buffer_avalon_pixel_dma_master_waitrequest   => pixel_buffer_avalon_pixel_dma_master_waitrequest,   --                                         .waitrequest
			pixel_buffer_avalon_pixel_dma_master_read          => pixel_buffer_avalon_pixel_dma_master_read,          --                                         .read
			pixel_buffer_avalon_pixel_dma_master_readdata      => pixel_buffer_avalon_pixel_dma_master_readdata,      --                                         .readdata
			pixel_buffer_avalon_pixel_dma_master_readdatavalid => pixel_buffer_avalon_pixel_dma_master_readdatavalid, --                                         .readdatavalid
			pixel_buffer_avalon_pixel_dma_master_lock          => pixel_buffer_avalon_pixel_dma_master_lock,          --                                         .lock
			onchip_mem_s1_address                              => mm_interconnect_0_onchip_mem_s1_address,            --                            onchip_mem_s1.address
			onchip_mem_s1_write                                => mm_interconnect_0_onchip_mem_s1_write,              --                                         .write
			onchip_mem_s1_readdata                             => mm_interconnect_0_onchip_mem_s1_readdata,           --                                         .readdata
			onchip_mem_s1_writedata                            => mm_interconnect_0_onchip_mem_s1_writedata,          --                                         .writedata
			onchip_mem_s1_byteenable                           => mm_interconnect_0_onchip_mem_s1_byteenable,         --                                         .byteenable
			onchip_mem_s1_chipselect                           => mm_interconnect_0_onchip_mem_s1_chipselect,         --                                         .chipselect
			onchip_mem_s1_clken                                => mm_interconnect_0_onchip_mem_s1_clken               --                                         .clken
		);

	mm_interconnect_1 : component lab2q_mm_interconnect_1
		port map (
			sys_sdram_pll_sys_clk_clk                             => sys_sdram_pll_sys_clk_clk,                                               --                      sys_sdram_pll_sys_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                                          --          cpu_reset_n_reset_bridge_in_reset.reset
			sysid_reset_reset_bridge_in_reset_reset               => rst_controller_002_reset_out_reset,                                      --          sysid_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                               => cpu_data_master_address,                                                 --                            cpu_data_master.address
			cpu_data_master_waitrequest                           => cpu_data_master_waitrequest,                                             --                                           .waitrequest
			cpu_data_master_byteenable                            => cpu_data_master_byteenable,                                              --                                           .byteenable
			cpu_data_master_read                                  => cpu_data_master_read,                                                    --                                           .read
			cpu_data_master_readdata                              => cpu_data_master_readdata,                                                --                                           .readdata
			cpu_data_master_write                                 => cpu_data_master_write,                                                   --                                           .write
			cpu_data_master_writedata                             => cpu_data_master_writedata,                                               --                                           .writedata
			cpu_data_master_debugaccess                           => cpu_data_master_debugaccess,                                             --                                           .debugaccess
			cpu_instruction_master_address                        => cpu_instruction_master_address,                                          --                     cpu_instruction_master.address
			cpu_instruction_master_waitrequest                    => cpu_instruction_master_waitrequest,                                      --                                           .waitrequest
			cpu_instruction_master_read                           => cpu_instruction_master_read,                                             --                                           .read
			cpu_instruction_master_readdata                       => cpu_instruction_master_readdata,                                         --                                           .readdata
			cpu_instruction_master_readdatavalid                  => cpu_instruction_master_readdatavalid,                                    --                                           .readdatavalid
			character_buffer_avalon_char_buffer_slave_address     => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_address,     --  character_buffer_avalon_char_buffer_slave.address
			character_buffer_avalon_char_buffer_slave_write       => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_write,       --                                           .write
			character_buffer_avalon_char_buffer_slave_read        => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_read,        --                                           .read
			character_buffer_avalon_char_buffer_slave_readdata    => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_readdata,    --                                           .readdata
			character_buffer_avalon_char_buffer_slave_writedata   => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_writedata,   --                                           .writedata
			character_buffer_avalon_char_buffer_slave_byteenable  => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_byteenable,  --                                           .byteenable
			character_buffer_avalon_char_buffer_slave_waitrequest => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_waitrequest, --                                           .waitrequest
			character_buffer_avalon_char_buffer_slave_chipselect  => mm_interconnect_1_character_buffer_avalon_char_buffer_slave_chipselect,  --                                           .chipselect
			character_buffer_avalon_char_control_slave_address    => mm_interconnect_1_character_buffer_avalon_char_control_slave_address,    -- character_buffer_avalon_char_control_slave.address
			character_buffer_avalon_char_control_slave_write      => mm_interconnect_1_character_buffer_avalon_char_control_slave_write,      --                                           .write
			character_buffer_avalon_char_control_slave_read       => mm_interconnect_1_character_buffer_avalon_char_control_slave_read,       --                                           .read
			character_buffer_avalon_char_control_slave_readdata   => mm_interconnect_1_character_buffer_avalon_char_control_slave_readdata,   --                                           .readdata
			character_buffer_avalon_char_control_slave_writedata  => mm_interconnect_1_character_buffer_avalon_char_control_slave_writedata,  --                                           .writedata
			character_buffer_avalon_char_control_slave_byteenable => mm_interconnect_1_character_buffer_avalon_char_control_slave_byteenable, --                                           .byteenable
			character_buffer_avalon_char_control_slave_chipselect => mm_interconnect_1_character_buffer_avalon_char_control_slave_chipselect, --                                           .chipselect
			cpu_jtag_debug_module_address                         => mm_interconnect_1_cpu_jtag_debug_module_address,                         --                      cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write                           => mm_interconnect_1_cpu_jtag_debug_module_write,                           --                                           .write
			cpu_jtag_debug_module_read                            => mm_interconnect_1_cpu_jtag_debug_module_read,                            --                                           .read
			cpu_jtag_debug_module_readdata                        => mm_interconnect_1_cpu_jtag_debug_module_readdata,                        --                                           .readdata
			cpu_jtag_debug_module_writedata                       => mm_interconnect_1_cpu_jtag_debug_module_writedata,                       --                                           .writedata
			cpu_jtag_debug_module_byteenable                      => mm_interconnect_1_cpu_jtag_debug_module_byteenable,                      --                                           .byteenable
			cpu_jtag_debug_module_waitrequest                     => mm_interconnect_1_cpu_jtag_debug_module_waitrequest,                     --                                           .waitrequest
			cpu_jtag_debug_module_debugaccess                     => mm_interconnect_1_cpu_jtag_debug_module_debugaccess,                     --                                           .debugaccess
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,                   --                jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,                     --                                           .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,                      --                                           .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,                  --                                           .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,                 --                                           .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,               --                                           .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,                --                                           .chipselect
			mouse_0_avalon_ps2_slave_address                      => mm_interconnect_1_mouse_0_avalon_ps2_slave_address,                      --                   mouse_0_avalon_ps2_slave.address
			mouse_0_avalon_ps2_slave_write                        => mm_interconnect_1_mouse_0_avalon_ps2_slave_write,                        --                                           .write
			mouse_0_avalon_ps2_slave_read                         => mm_interconnect_1_mouse_0_avalon_ps2_slave_read,                         --                                           .read
			mouse_0_avalon_ps2_slave_readdata                     => mm_interconnect_1_mouse_0_avalon_ps2_slave_readdata,                     --                                           .readdata
			mouse_0_avalon_ps2_slave_writedata                    => mm_interconnect_1_mouse_0_avalon_ps2_slave_writedata,                    --                                           .writedata
			mouse_0_avalon_ps2_slave_byteenable                   => mm_interconnect_1_mouse_0_avalon_ps2_slave_byteenable,                   --                                           .byteenable
			mouse_0_avalon_ps2_slave_waitrequest                  => mm_interconnect_1_mouse_0_avalon_ps2_slave_waitrequest,                  --                                           .waitrequest
			mouse_0_avalon_ps2_slave_chipselect                   => mm_interconnect_1_mouse_0_avalon_ps2_slave_chipselect,                   --                                           .chipselect
			pixel_buffer_avalon_control_slave_address             => mm_interconnect_1_pixel_buffer_avalon_control_slave_address,             --          pixel_buffer_avalon_control_slave.address
			pixel_buffer_avalon_control_slave_write               => mm_interconnect_1_pixel_buffer_avalon_control_slave_write,               --                                           .write
			pixel_buffer_avalon_control_slave_read                => mm_interconnect_1_pixel_buffer_avalon_control_slave_read,                --                                           .read
			pixel_buffer_avalon_control_slave_readdata            => mm_interconnect_1_pixel_buffer_avalon_control_slave_readdata,            --                                           .readdata
			pixel_buffer_avalon_control_slave_writedata           => mm_interconnect_1_pixel_buffer_avalon_control_slave_writedata,           --                                           .writedata
			pixel_buffer_avalon_control_slave_byteenable          => mm_interconnect_1_pixel_buffer_avalon_control_slave_byteenable,          --                                           .byteenable
			sdram_controller_s1_address                           => mm_interconnect_1_sdram_controller_s1_address,                           --                        sdram_controller_s1.address
			sdram_controller_s1_write                             => mm_interconnect_1_sdram_controller_s1_write,                             --                                           .write
			sdram_controller_s1_read                              => mm_interconnect_1_sdram_controller_s1_read,                              --                                           .read
			sdram_controller_s1_readdata                          => mm_interconnect_1_sdram_controller_s1_readdata,                          --                                           .readdata
			sdram_controller_s1_writedata                         => mm_interconnect_1_sdram_controller_s1_writedata,                         --                                           .writedata
			sdram_controller_s1_byteenable                        => mm_interconnect_1_sdram_controller_s1_byteenable,                        --                                           .byteenable
			sdram_controller_s1_readdatavalid                     => mm_interconnect_1_sdram_controller_s1_readdatavalid,                     --                                           .readdatavalid
			sdram_controller_s1_waitrequest                       => mm_interconnect_1_sdram_controller_s1_waitrequest,                       --                                           .waitrequest
			sdram_controller_s1_chipselect                        => mm_interconnect_1_sdram_controller_s1_chipselect,                        --                                           .chipselect
			sysid_control_slave_address                           => mm_interconnect_1_sysid_control_slave_address,                           --                        sysid_control_slave.address
			sysid_control_slave_readdata                          => mm_interconnect_1_sysid_control_slave_readdata                           --                                           .readdata
		);

	irq_mapper : component lab2q_irq_mapper
		port map (
			clk           => sys_sdram_pll_sys_clk_clk,      --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component lab2q_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_reset_source_reset,   -- reset_in0.reset
			clk            => sys_sdram_pll_sys_clk_clk,          --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component lab2q_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => video_clk_reset_source_reset,       -- reset_in0.reset
			clk            => video_clk_vga_clk_clk,              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component lab2q_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => sys_sdram_pll_sys_clk_clk,          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_1_sdram_controller_s1_read_ports_inv <= not mm_interconnect_1_sdram_controller_s1_read;

	mm_interconnect_1_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_1_sdram_controller_s1_byteenable;

	mm_interconnect_1_sdram_controller_s1_write_ports_inv <= not mm_interconnect_1_sdram_controller_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of lab2q
